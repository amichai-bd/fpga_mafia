//------------------------------------
// Project:   CPUC
// File name: cpuc.sv
// Date:      26.12.24
// Author:     
//--------------------------------------
// Description: cpuc grid
//--------------------------------------

`include "cpuc_macros.vh"

module cpuc 
import cpuc_package::*;
(
    input logic clk,
    input logic rst,
    output var t_reg_outputs reg_output
);



endmodule