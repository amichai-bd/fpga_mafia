module cpuc_tb;

initial begin
    #10
    $finish;
end

endmodule